library verilog;
use verilog.vl_types.all;
entity bcd_3digit_incrementor_tb is
end bcd_3digit_incrementor_tb;
