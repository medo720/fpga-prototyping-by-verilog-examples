library verilog;
use verilog.vl_types.all;
entity sign_mag_add_test is
end sign_mag_add_test;
