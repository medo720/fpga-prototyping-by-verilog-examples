library verilog;
use verilog.vl_types.all;
entity eq1 is
    port(
        i0              : in     vl_logic;
        i1              : in     vl_logic;
        eq              : out    vl_logic
    );
end eq1;
