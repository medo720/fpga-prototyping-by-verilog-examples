library verilog;
use verilog.vl_types.all;
entity eq2_testbench is
end eq2_testbench;
